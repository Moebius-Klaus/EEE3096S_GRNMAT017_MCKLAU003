`timescale 1ns / 1ps

module alu( clk, operand_a, operand_b, opcode, result);
    parameter DATA_WIDTH = 8;

    input clk;
    input[DATA_WIDTH-1:0]operand_a,operand_b;
    input [3:0] opcode;
    output reg[DATA_WIDTH-1:0] result;
    
  always@(posedge clk)
    begin
     case(opcode)
        4'b0000: //Addition
           result <= operand_a + operand_b ; 
        4'b0001: //Subtraction 
           result <= operand_a - operand_b;
        default: result <= 8'bx; 
     endcase
     
    end
endmodule